module statistic( clock, reset, clear, DataIn1, DataIn2, EvenParity, GreyCode, overflow);
input clock; // Clock
input reset; // synchronous reset - active low
input clear; // Clears statistics when high (synchronous)
input [7:0] DataIn1; // Input Data 1
input [7:0] DataIn2; // Input Data 2
// all outputs are registered 
output [7:0] EvenParity; // # of data with Even parity 
output [7:0] GreyCode; // # of data with pattern 10101010 or 01010101    
output overflow; // =1 if any of the counters above overflow, stays high until clear goes high
reg [7:0] GreyCode, EvenParity;
reg overflow;
wire In1, In2;
reg Grey1, Grey2;
wire adder_carry_1, adder_carry_2;
wire [7:0] Sum1, Sum2;

always@(posedge clock) 
begin

if(!reset)
begin
GreyCode<=0;
EvenParity <= 0;
overflow <=0;
end 

else if(clear)
begin
GreyCode<=0;
EvenParity <= 0;
overflow <=0;
end 

else
begin
overflow <= (overflow | (adder_carry_1 | adder_carry_2));
EvenParity <= Sum1;
GreyCode <= Sum2;
end 
end

assign In1 = ~(^DataIn1);
assign In2 = ~(^DataIn2);

assign{ adder_carry_1,Sum1} = In1+In2+ EvenParity;
assign{ adder_carry_2,Sum2} = Grey1+Grey2+GreyCode;

always@(*)
begin
Grey1 = 0; Grey2 = 0; 
if((DataIn1==8'b10101010)||(DataIn1==8'b01010101))
Grey1 = 1;
if((DataIn2==8'b01010101)||(DataIn2==8'b10101010))
Grey2 = 1;
end

endmodule

